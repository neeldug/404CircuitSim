* D:\home\jjl119\Imperial\SummerProject\404CircuitSim\test\SpiceNetlists\Draft4.asc
V1 N001 N003 SINE(0 10 1000)
R1 N002 0 1000
D1 0 N001 D
D2 N001 N002 D
D3 0 N003 D
D4 N003 N002 D
C1 N002 0 1n
.model D D
.lib C:\users\jjl119\My Documents\LTspiceXVII\lib\cmp\standard.dio
.tran 0 3m 0 0.001m
.backanno
.end
