* D:\home\jjl119\Imperial\SummerProject\404CircuitSim\test\SpiceNetlists\Draft4.asc
V1 N001 0 SINE(0 5 1000)
R2 N002 N001 1000
D1 N002 0 D
.tran 0 1m 0 0.01m
.backanno
.end
