* Voltage Sources
V1 N001 0 5
R1 N002 N001 10
R2 N003 N002 1k
C1 N002 0 0.1m
L1 N003 0 100m
.tran 0 1 0 0.1m
.backanno
.end
