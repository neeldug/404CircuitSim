* D:\home\jjl119\Imperial\SummerProject\404CircuitSim\test\SpiceNetlists\Draft4.asc
V1 N001 0 SINE(0 5 1000)
D1 N001 N002 D
R1 N002 0 1000
C1 N002 0 1n
.model D D
.lib C:\users\jjl119\My Documents\LTspiceXVII\lib\cmp\standard.dio
.tran 0 1m 0 0.01m
.backanno
.end
