D:\home\jjl119\Imperial\SummerProject\404CircuitSim\test\SpiceNetlists\Draft4.asc
V1 N001 0 5
R2 N002 N001 10
C1 N002 0 10u
.tran 0 10m 0 0.005m
.backanno
.end
