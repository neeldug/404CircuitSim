*Title
C1 N001 0 1u
R1 N001 0 100000
I1 N001 0 50u
.tran 0 1 0 1u
.backanno
.end