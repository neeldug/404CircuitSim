* D:\home\jjl119\Imperial\SummerProject\404CircuitSim\test\SpiceNetlists\Draft4.asc
R1 N001 0 {R}
V1 N001 0 SINE(0 1 1000)
.step param R 1 10 1
.tran 0 2m 0 0.01m
.backanno
.end
