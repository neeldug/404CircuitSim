* D:\home\jjl119\Imperial\SummerProject\404CircuitSim\test\SpiceNetlists\Draft4.asc
D1 0 N001 D
D2 0 N003 D
D4 N003 N002 D
R1 N002 0 {R}
V2 N001 N003 SINE(0 5 1000)
D3 N001 N002 D
.model D D
.step DEC param R 10 10000 1
.tran 0 10m 0 0.01m
.backanno
.end
