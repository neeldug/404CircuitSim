* C:\users\sam\My Documents\LTspiceXVII\Draft1.asc
R1 N003 0 1
V1 N001 0 SINE(0 5 1k)
R2 N003 N001 1
R3 N002 N001 1
R4 N002 N003 1
R5 N003 N002 1
V2 N003 N004 5
R6 N004 0 1
.tran 0 0.2 0 0.01m
.backanno
.end
