* D:\home\jjl119\Imperial\SummerProject\404CircuitSim\Draft1.asc
V1 N001 N002 5
R1 N001 N002 5
.backanno
.end

