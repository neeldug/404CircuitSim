* D:\home\jjl119\Imperial\SummerProject\404CircuitSim\test\SpiceNetlists\Draft4.asc
R1 N002 N001 1000
C1 N002 0 10n
V1 N001 0 5
.tran 0 10u 0 0.01u
.backanno
.end
