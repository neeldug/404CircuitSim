*50
V1 1 0 SINE(0 100 1)
R1 1 2 1
R51 1 0 1000
R2 2 3 1
R52 2 0 1000
R3 3 4 1
R53 3 0 1000
R4 4 5 1
R54 4 0 1000
R5 5 6 1
R55 5 0 1000
R6 6 7 1
R56 6 0 1000
R7 7 8 1
R57 7 0 1000
R8 8 9 1
R58 8 0 1000
R9 9 10 1
R59 9 0 1000
R10 10 11 1
R60 10 0 1000
R11 11 12 1
R61 11 0 1000
R12 12 13 1
R62 12 0 1000
R13 13 14 1
R63 13 0 1000
R14 14 15 1
R64 14 0 1000
R15 15 16 1
R65 15 0 1000
R16 16 17 1
R66 16 0 1000
R17 17 18 1
R67 17 0 1000
R18 18 19 1
R68 18 0 1000
R19 19 20 1
R69 19 0 1000
R20 20 21 1
R70 20 0 1000
R21 21 22 1
R71 21 0 1000
R22 22 23 1
R72 22 0 1000
R23 23 24 1
R73 23 0 1000
R24 24 25 1
R74 24 0 1000
R25 25 26 1
R75 25 0 1000
R26 26 27 1
R76 26 0 1000
R27 27 28 1
R77 27 0 1000
R28 28 29 1
R78 28 0 1000
R29 29 30 1
R79 29 0 1000
R30 30 31 1
R80 30 0 1000
R31 31 32 1
R81 31 0 1000
R32 32 33 1
R82 32 0 1000
R33 33 34 1
R83 33 0 1000
R34 34 35 1
R84 34 0 1000
R35 35 36 1
R85 35 0 1000
R36 36 37 1
R86 36 0 1000
R37 37 38 1
R87 37 0 1000
R38 38 39 1
R88 38 0 1000
R39 39 40 1
R89 39 0 1000
R40 40 41 1
R90 40 0 1000
R41 41 42 1
R91 41 0 1000
R42 42 43 1
R92 42 0 1000
R43 43 44 1
R93 43 0 1000
R44 44 45 1
R94 44 0 1000
R45 45 46 1
R95 45 0 1000
R46 46 47 1
R96 46 0 1000
R47 47 48 1
R97 47 0 1000
R48 48 49 1
R98 48 0 1000
R49 49 50 1
R99 49 0 1000
.tran 0 3 0 0.001
.end
