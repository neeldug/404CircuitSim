* C:\users\jjl119\My Documents\LTspiceXVII\Draft2.asc
R1 N001 N003 1000
R2 N001 N002 2000
C1 N003 0 10n
L1 N002 0 1m
I1 0 N001 SINE(0 1m 1000)
.tran 0 50m 2m 0.01m
.backanno
.end
