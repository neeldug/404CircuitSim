* C:\users\jjl119\My Documents\LTspiceXVII\Draft1.asc
V1 N001 N002 SINE(1 4 2)
R1 N001 N002 10
.backanno
.end

