* C:\users\jjl119\My Documents\LTspiceXVII\Draft1.asc
V1 N001 N004 1
V2 N002 N004 AC 2
V3 N003 N004 SINE(3 4 5)
R1 0 N001 1000
L1 0 N002 2000
C1 0 N003 3000
I1 N004 N005 6
I2 N004 N006 AC 7
I3 N004 N007 SINE(8 9 10)
R2 N005 0 4000
R3 N006 0 5000
R4 N007 0 6000
.backanno
.end
