* D:\home\jjl119\Imperial\SummerProject\404CircuitSim\test\SpiceNetlists\Draft4.asc
V1 N001 0 SINE(0 10 1000)
R1 N002 0 1000
D1 N001 N002 D
D2 N002 N001 D
.model D D
.tran 0 3m 0 0.01m
.backanno
.end
